library ieee;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity memory is
  port (
    dir : in std_logic_vector (11 downto 0);
    data : out std_logic_vector (93 downto 0));

end memory;

architecture behavioral of memory is

begin
  process(dir)
  begin

    -- data format
    -- |    prueba    |vf| ins |                liga                 |
    --  p4 p3 p2 p1 p0 vf i1 i0 l11 l10 l9 l8 l7 l6 l5 l4 l3 l2 l1 l0 ncri eb1 eb0 nwb ea1 ea0 nwa selbus upa9 upa8 upa7 upa6 upa5 upa4 upa3 upa2 upa1 upa0 noeupa ndupa selmux nex2 nex1 nex0 x2 x1 x0 enay nera2 nera1 nera0 ra2 ra1 ra0 neap2 neap1 neap0 ap2 ap1 ap0 nepc2 nepc1 nepc0 pc2 pc1 pc0 ncbd nas nrw bd dint hint set_irq set_xirq b9 b8 b7 b6 b5 b4 b3 b2 b1 b0 cc cn cv cz ci ch cx cs nhb accsec
	--ciclo fetch
    case dir is
      when x"000" => data <= "0000000000000000000010010010000000000011011100001110001110000110000110000000000000000000000010";
      when x"001" => data <= "0000000000000000000000010010000000000011011100001110001110001110011010000000000000000000000010";
      when x"002" => data <= "0000001000000000000010010010000000000011011100001110001110001110001110000000000000000000000010";

      -- cba (acceso inherente) n,z,v,c
      when x"110" => data <= "0000000000000000000011111110001010000111111100001110001110001110001110000000000000000000000011";
      -- eb1,eb0,ea1,ea0,upa7,upa5,upa0,selmux,accsec
      when x"111" => data <= "0000000000000000000010010010000000000000011100001110001110001110001110000000000000000000000010";
      when x"112" => data <= "0111111100000000000010010010000000000011011100001110001110001110001110000000000000001111000010";
      -- cc,cv,cn,cz,salto de interrupción (mi=11, prueba=15 int)
      when x"113" => data <= "1100000100000000000110010010000000000011011100001110001110000110000110000000000000000000000010";
		     -- salto condicional (mi=01, prueba=24 0), salto a x"001", nepc2,ncbd

      -- ja (acceso directo)
      when x"270" => data <= "0000000000000000000010011110000100000011011100001110001110001110001110000000000000000000000010";
      -- upa6,ea0,ea1
      when x"271" => data <= "0000000000000000000010010010000000000000011100001011001110001110001110000000000000000000000010";
      -- ra2,nera1,ndupa,noeupa
      when x"272" => data <= "0000000000000000000010010010000000000011011100001110001110000110000110000000000000000000000010";
      -- nepc2,ncbd
      when x"273" => data <= "0000000000000000000010010010000000000011011100001100111110001110001010000000000000000000000010";
      -- nas,nera0,ra1,ra0
      when x"274" => data <= "0000000000000000000010010010000000000011011100000110001110001110010110000000000000000000000010";
      -- nera2,ncbd,pc0
      when x"275" => data <= "1000000100100111011110010010000000000011011100001110001110001110001110000000000000000000000010";
      -- salto condicional (mi=01, prueba=16 c) salto a x"277"=001001110111
      when x"276" => data <= "0000000000000000000010010010000000000011011100001000001110001001011110000000000000000000000010";
      -- nepc1,nepc0,nera1,nera0,pc2,pc0
      when x"277" => data <= "1100000100000000000110010010000000000011011100001110001110000110000110000000000000000000000010";
		     -- salto condicional (mi=01, prueba=24 0), salto a x"001", nepc2,ncbd

      -- staa (acceso directo)
      when x"970" => data <= "0000000000000000000010011110000100000011011100001110001110001110001110000000000000000000000010";
      -- upa6,ea0,ea1
      when x"971" => data <= "0000000000000000000010010010000000000000011100001011001110001110001110000000000000000000000010";
      -- ra2,nera1,ndupa,noeupa
      when x"972" => data <= "0000000000000000000010010010000000000011011100001110001110000110000110000000000000000000000010";
      -- nepc2,ncbd
      when x"973" => data <= "0000000000000000000010010010000000000011011100001100111110001110001010000000000000000000000010";
      -- nas,nera0,ra1,ra0
      when x"974" => data <= "0000000000000000000010010010000000000011011100000110001110001110010110000000000000000000000010";
      -- nera2,ncbd,pc0
      when x"975" => data <= "0000000000000000000010010110000000000011011100001110001110001110001000000000000000000000000010";
      -- nrw,nas,ea0
      when x"976" => data <= "0000000000000000000010010010000000000011011100001110001110001110001110000000010011000000000010";
      when x"977" => data <= "0111111100000000000010010010000000000011011100001110001110001110001110000000010011000111000010";
      -- b6,b3,b2,cn,cv,cz,salto de interrupción (mi=11, prueba=15 int)
      when x"978" => data <= "1100000100000000000110010010000000000011011100001110001110000110000110000000000000000000000010";
		     -- salto condicional (mi=01, prueba=24 0), salto a x"001", nepc2,ncbd

      -- stab (acceso directo)
      when x"d70" => data <= "0000000000000000000010011110000100000011011100001110001110001110001110000000000000000000000010";
      -- upa6,ea0,ea1
      when x"d71" => data <= "0000000000000000000010010010000000000000011100001011001110001110001110000000000000000000000010";
      -- ra2,nera1,ndupa,noeupa
      when x"d72" => data <= "0000000000000000000010010010000000000011011100001110001110000110000110000000000000000000000010";
      -- nepc2,ncbd
      when x"d73" => data <= "0000000000000000000010010010000000000011011100001100111110001110001010000000000000000000000010";
      -- nas,nera0,ra1,ra0
      when x"d74" => data <= "0000000000000000000010010010000000000011011100000110001110001110010110000000000000000000000010";
      -- nera2,ncbd,pc0
      when x"d75" => data <= "0000000000000000000010110010000000000011011100001110001110001110001000000000000000000000000010";
      -- nrw,nas,eb0
      when x"d77" => data <= "0111111100000000000010010010000000000011011100001110001110001110001110000000100101000111000010";
      -- b7,b4,b2,cn,cv,cz,salto de interrupción (mi=11, prueba=15 int)
      when x"d78" => data <= "1100000100000000000110010010000000000011011100001110001110000110000110000000000000000000000010";
		     -- salto condicional (mi=01, prueba=24 0), salto a x"001", nepc2,ncbd

      -- ldaa (acceso directo)
      when x"960" => data <= "0000000000000000000010011110000100000011011100001110001110001110001110000000000000000000000010";
      -- upa6,ea0,ea1
      when x"961" => data <= "0000000000000000000010010010000000000000011100001011001110001110001110000000000000000000000010";
      -- ra2,nera1,ndupa,noeupa
      when x"962" => data <= "0000000000000000000010010010000000000011011100001110001110000110000110000000000000000000000010";
      -- nepc2,ncbd
      when x"963" => data <= "0000000000000000000010010010000000000011011100001100111110001110001010000000000000000000000010";
      -- nas,nera0,ra1,ra0
      when x"964" => data <= "0000000000000000000010010010000000000011011100000110001110001110010110000000000000000000000010";
      -- nera2,ncbd.pc0
      when x"965" => data <= "0000000000000000000010010100000000000011011100001110001110001110001010000000000000000000000010";
      -- nas,ea0,nwa
      when x"967" => data <= "0111111100000000000010010010000000000011011100001110001110001110001110000000010011000111000010";
      -- b6,b3,b2,cn,cv,cz,salto de interrupción (mi=11, prueba=15 int)
      when x"968" => data <= "1100000100000000000110010010000000000011011100001110001110000110000110000000000000000000000010";
		     -- salto condicional (mi=01, prueba=24 0), salto a x"001", nepc2,ncbd


      --ldaa(acceso inmediato)
      when x"860" => data <= "0000000000000000000010010010000000000011011100001110001110000110000110000000000000000000000010";
      when x"861" => data <= "0000000000000000000010010100000000000011011100001110001110001110011010000000000000000000000010";
      when x"862" => data <= "0111111100000000000010010010000000000011011100001110001110001110001110000000010011000111000010";
      when x"863" => data <= "1100000100000000000110010010000000000011011100001110001110000110000110000000000000000000000010";

      -- ldab (acceso directo)
      when x"d60" => data <= "0000000000000000000010011110000100000011011100001110001110001110001110000000000000000000000010";
      -- upa6,ea0,ea1
      when x"d61" => data <= "0000000000000000000010010010000000000000011100001011001110001110001110000000000000000000000010";
      -- ra2,nera1,ndupa,noeupa
      when x"d62" => data <= "0000000000000000000010010010000000000011011100001110001110000110000110000000000000000000000010";
      -- nepc2,ncbd
      when x"d63" => data <= "0000000000000000000010010010000000000011011100001100111110001110001010000000000000000000000010";
      -- nas,nera0,ra1,ra0
      when x"d64" => data <= "0000000000000000000010010010000000000011011100000110001110001110010110000000000000000000000010";
      -- nera2,ncbd,pc0
      when x"d65" => data <= "0000000000000000000010100010000000000011011100001110001110001110001010000000000000000000000010";
      -- nas,eb0,nwb
      when x"d67" => data <= "0111111100000000000010010010000000000011011100001110001110001110001110000000100101000111000010";
      -- b7,b4,b2,cn,cv,cz,salto de interrupción (mi=11, prueba=15 int)
      when x"d68" => data <= "1100000100000000000110010010000000000011011100001110001110000110000110000000000000000000000010";
		     -- salto condicional (mi=01, prueba=24 0), salto a x"001", nepc2,ncbd


      --ldab(acceso inmediato)
      when x"c60" => data <= "0000000000000000000010010010000000000011011100001110001110000110000110000000000000000000000010";
      when x"c61" => data <= "0000000000000000000010100010000000000011011100001110001110001110011010000000000000000000000010";
      when x"c62" => data <= "0111111100000000000010010010000000000011011100001110001110001110001110000000100101000111000010";
      when x"c63" => data <= "1100000100000000000110010010000000000011011100001110001110000110000110000000000000000000000010";

      -- aba a=a+b (inherente)
      when x"1b0" => data <= "0000000000000000000011111110000000000111111100001110001110001110001110000000000000000000000010";
      when x"1b1" => data <= "0111111100000000000010010100000000000000011100001110001110001110001110000000000000001111010010";
      when x"1b2" => data <= "1100000100000000000110010010000000000011011100001110001110000110000110000000000000000000000010";

      --jum acceso (ext)
      when x"7e0" => data <= "0000000000000000000010010010000000000011011100001110001110000110000110000000000000000000000010";
      when x"7e1" => data <= "0000000000000000000010010010000000000011011100001011001110001110011011000000000000000000000010";
      when x"7e2" => data <= "0000000000000000000010010010000000000011011100001110001110000110000110000000000000000000000010";
      when x"7e3" => data <= "0000000000000000000010010010000000000011011100001100111110001110011010000000000000000000000010";
      when x"7e4" => data <= "0111111100000000000010010010000000000011011100001000001110001001011110000000000000000000000010";
      when x"7e5" => data <= "1100000100000000000110010010000000000011011100001110001110000110000110000000000000000000000010";

		when others => data <= "0000000000000000000010010010000000000011011100001110001110001110001110000000000000000000000010";
		 -- default

    end case;

  end process;
end behavioral;
